module mux4to1_case (
    input  wire [1:0] sel,
    input  wire [3:0] in,
    output reg        out
);
    always @(*) begin
        case (sel)
            2'b00: out = in[0];
            2'b01: out = in[1];
            2'b10: out = in[2];
            2'b11: out = in[3];
        endcase
    end
endmodule